<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-130.333,-521.211,64.0667,-619.477</PageViewport>
<gate>
<ID>389</ID>
<type>AA_TOGGLE</type>
<position>-101,-426</position>
<output>
<ID>OUT_0</ID>219 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>390</ID>
<type>AA_TOGGLE</type>
<position>-87,-426</position>
<output>
<ID>OUT_0</ID>220 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>391</ID>
<type>AA_LABEL</type>
<position>-93.5,-418.5</position>
<gparam>LABEL_TEXT 1.Using AOI gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>392</ID>
<type>AA_INVERTER</type>
<position>-95.5,-429.5</position>
<input>
<ID>IN_0</ID>219 </input>
<output>
<ID>OUT_0</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>393</ID>
<type>AA_INVERTER</type>
<position>-82.5,-430.5</position>
<input>
<ID>IN_0</ID>220 </input>
<output>
<ID>OUT_0</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_LABEL</type>
<position>-101,-423</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>395</ID>
<type>AA_LABEL</type>
<position>-87,-423</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>AA_AND2</type>
<position>-60.5,-437</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_AND2</type>
<position>-60,-446.5</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>AE_OR2</type>
<position>-50,-440.5</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>GA_LED</type>
<position>-42.5,-440.5</position>
<input>
<ID>N_in0</ID>225 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>-28.5,-439.5</position>
<gparam>LABEL_TEXT D=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>AA_LABEL</type>
<position>-30.5,-436.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>AA_LABEL</type>
<position>-22,-436.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>GA_LED</type>
<position>-42,-454.5</position>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>AA_LABEL</type>
<position>-32,-454</position>
<gparam>LABEL_TEXT Bo=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>407</ID>
<type>AA_AND2</type>
<position>-58,-455</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_LABEL</type>
<position>-30,-451</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>409</ID>
<type>AA_LABEL</type>
<position>6.5,-419</position>
<gparam>LABEL_TEXT 2.Using NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>AA_TOGGLE</type>
<position>-5,-427</position>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_TOGGLE</type>
<position>8.5,-427</position>
<output>
<ID>OUT_0</ID>228 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>8,6.5</position>
<gparam>LABEL_TEXT Basic logic gates</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>412</ID>
<type>GA_LED</type>
<position>44.5,-438.5</position>
<input>
<ID>N_in0</ID>233 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>413</ID>
<type>AA_LABEL</type>
<position>56.5,-437.5</position>
<gparam>LABEL_TEXT D=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>414</ID>
<type>AA_LABEL</type>
<position>54.5,-434.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>415</ID>
<type>AA_LABEL</type>
<position>63,-434.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>416</ID>
<type>GA_LED</type>
<position>46,-453</position>
<input>
<ID>N_in2</ID>237 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>417</ID>
<type>AA_LABEL</type>
<position>55.5,-452.5</position>
<gparam>LABEL_TEXT Bo=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>-5,-424</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>419</ID>
<type>BA_NAND2</type>
<position>14,-431</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_LABEL</type>
<position>9,-424</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>-46,-8.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>BA_NAND2</type>
<position>1.5,-431.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-57,-6</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>422</ID>
<type>BA_NAND2</type>
<position>26.5,-436</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-57,-11</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>423</ID>
<type>BA_NAND2</type>
<position>27,-442.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>-38,-8</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>BA_NAND2</type>
<position>37,-438.5</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>-61.5,-5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>-61.5,-10.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>BA_NAND2</type>
<position>28,-453</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>428</ID>
<type>BA_NAND2</type>
<position>37.5,-453</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>AA_LABEL</type>
<position>57.5,-449.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>430</ID>
<type>AA_LABEL</type>
<position>-91,-465</position>
<gparam>LABEL_TEXT 3.Using NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>431</ID>
<type>AA_TOGGLE</type>
<position>-103.5,-475</position>
<output>
<ID>OUT_0</ID>238 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>432</ID>
<type>AA_TOGGLE</type>
<position>-86.5,-475</position>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>433</ID>
<type>GA_LED</type>
<position>-44.5,-488</position>
<input>
<ID>N_in1</ID>245 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>-60.5,-1.5</position>
<gparam>LABEL_TEXT 1.AND gates</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>-34.5,-484.5</position>
<gparam>LABEL_TEXT D=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>-36.5,-481.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>AA_LABEL</type>
<position>-28,-481.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>GA_LED</type>
<position>-50.5,-501</position>
<input>
<ID>N_in2</ID>247 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>438</ID>
<type>AA_LABEL</type>
<position>-41.5,-500.5</position>
<gparam>LABEL_TEXT Bo=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>-104,-472</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>-86.5,-472</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>441</ID>
<type>BE_NOR2</type>
<position>-97.5,-480</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>442</ID>
<type>BE_NOR2</type>
<position>-79.5,-478.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>BE_NOR2</type>
<position>-69,-484.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>444</ID>
<type>BE_NOR2</type>
<position>-68.5,-492.5</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>445</ID>
<type>BE_NOR2</type>
<position>-59.5,-488</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>446</ID>
<type>BE_NOR2</type>
<position>-50.5,-488</position>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>448</ID>
<type>AA_LABEL</type>
<position>-39.5,-497</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>449</ID>
<type>BE_NOR2</type>
<position>-68,-501</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>451</ID>
<type>AA_LABEL</type>
<position>-40,-515.5</position>
<gparam>LABEL_TEXT FULL ADDER</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>452</ID>
<type>AA_TOGGLE</type>
<position>-95,-533</position>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_TOGGLE</type>
<position>-80.5,-533</position>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>-58,-24</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>454</ID>
<type>AA_LABEL</type>
<position>-88,-525.5</position>
<gparam>LABEL_TEXT 1.Using AOI gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>-58,-29</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>-95.5,-530</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>-37.5,-26</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>-80.5,-529.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>-62,-23.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>457</ID>
<type>AA_TOGGLE</type>
<position>-64.5,-533.5</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>-62,-28.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AA_LABEL</type>
<position>-65,-530</position>
<gparam>LABEL_TEXT Cin</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>-61,-19</position>
<gparam>LABEL_TEXT 2.OR gates</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>-28,-7.5</position>
<gparam>LABEL_TEXT Y=A.B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>-28.5,-25.5</position>
<gparam>LABEL_TEXT Y=A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>462</ID>
<type>AE_SMALL_INVERTER</type>
<position>-91.5,-536</position>
<input>
<ID>IN_0</ID>248 </input>
<output>
<ID>OUT_0</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_SMALL_INVERTER</type>
<position>-76,-536</position>
<input>
<ID>IN_0</ID>249 </input>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_OR2</type>
<position>-46,-26</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>AE_SMALL_INVERTER</type>
<position>-59.5,-536.5</position>
<input>
<ID>IN_0</ID>250 </input>
<output>
<ID>OUT_0</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>-61,-58</position>
<gparam>LABEL_TEXT 4.XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>466</ID>
<type>AA_AND3</type>
<position>-49,-540</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>252 </input>
<input>
<ID>IN_2</ID>250 </input>
<output>
<ID>OUT</ID>258 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>467</ID>
<type>AA_AND3</type>
<position>-48.5,-550.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>253 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>468</ID>
<type>AA_AND3</type>
<position>-48,-560.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>252 </input>
<input>
<ID>IN_2</ID>253 </input>
<output>
<ID>OUT</ID>256 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_AND3</type>
<position>-47.5,-570</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>250 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>471</ID>
<type>AE_OR4</type>
<position>-29,-548.5</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>255 </input>
<input>
<ID>IN_2</ID>256 </input>
<input>
<ID>IN_3</ID>257 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>-59,-64.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>-59,-69</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>473</ID>
<type>GA_LED</type>
<position>-17.5,-548.5</position>
<input>
<ID>N_in0</ID>259 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>-37,-67</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>AA_LABEL</type>
<position>1.5,-545</position>
<gparam>LABEL_TEXT sum=ABCin+ABCin+ABCin+ABCin</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-63,-63.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>475</ID>
<type>AA_LABEL</type>
<position>-14.5,-542</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-63,-68.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>476</ID>
<type>AA_LABEL</type>
<position>-12.5,-542</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-26,-66.5</position>
<gparam>LABEL_TEXT Y=AB+BA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>477</ID>
<type>AA_LABEL</type>
<position>-3.5,-542</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>478</ID>
<type>AA_LABEL</type>
<position>0.5,-542</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>-62,-36</position>
<gparam>LABEL_TEXT 3.NOT gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>479</ID>
<type>AA_LABEL</type>
<position>9.5,-542</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>-58.5,-44.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_LABEL</type>
<position>12,-542</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>481</ID>
<type>AA_AND3</type>
<position>-47,-581.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>250 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_SMALL_INVERTER</type>
<position>-46,-44.5</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>-37,-44.5</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>483</ID>
<type>AA_AND3</type>
<position>-46.5,-600</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>253 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>-27,-43.5</position>
<gparam>LABEL_TEXT Y=A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>-62.5,-44</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>-25,-40.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>486</ID>
<type>AA_AND3</type>
<position>-46.5,-591.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>252 </input>
<input>
<ID>IN_2</ID>250 </input>
<output>
<ID>OUT</ID>262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>98</ID>
<type>AI_XOR2</type>
<position>-44.5,-67</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>488</ID>
<type>AE_OR4</type>
<position>-25,-588.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>262 </input>
<input>
<ID>IN_2</ID>263 </input>
<input>
<ID>IN_3</ID>266 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>-28,-63.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>489</ID>
<type>GA_LED</type>
<position>-14.5,-588.5</position>
<input>
<ID>N_in3</ID>265 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>-22,-63</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>490</ID>
<type>AA_LABEL</type>
<position>5.5,-584.5</position>
<gparam>LABEL_TEXT carry=ABCin+ABCin+ABCin+ABCin</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>8,-2.5</position>
<gparam>LABEL_TEXT 5.X-NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>491</ID>
<type>AA_LABEL</type>
<position>-10,-581.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>4.5,-8</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_LABEL</type>
<position>3.5,-581.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>4.5,-12.5</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>493</ID>
<type>AA_LABEL</type>
<position>17,-581.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>26.5,-10.5</position>
<input>
<ID>N_in3</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>0.5,-7</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>495</ID>
<type>AA_AND3</type>
<position>-46.5,-608.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<input>
<ID>IN_2</ID>250 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>0.5,-12</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>37.5,-10.5</position>
<gparam>LABEL_TEXT Y=AB+BA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>41.5,-7</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AO_XNOR2</type>
<position>17.5,-10</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>43.5,-7</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>-5,-84.5</position>
<gparam>LABEL_TEXT NAND gate as universal gate gate</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>-61,-99</position>
<gparam>LABEL_TEXT 1.NAND as NOT gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>BA_NAND2</type>
<position>-60.5,-107.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_TOGGLE</type>
<position>-70,-107.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>123</ID>
<type>GA_LED</type>
<position>-51.5,-108</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>-73,-107</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>-45.5,-107.5</position>
<gparam>LABEL_TEXT Y=A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>-43.5,-104.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-61.5,-115.5</position>
<gparam>LABEL_TEXT 2.NAND as AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>BA_NAND2</type>
<position>-60.5,-125</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>-70,-123</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>-42,-125</position>
<input>
<ID>N_in0</ID>59 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>-73,-122.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>-34,-124.5</position>
<gparam>LABEL_TEXT Y=A.B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>-69.5,-127.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>-73,-127</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>BA_NAND2</type>
<position>-50,-125</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>-63,-135</position>
<gparam>LABEL_TEXT 3.NAND as OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>BA_NAND2</type>
<position>-62,-144</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>-71,-144</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>-43.5,-144</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>-74,-143</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>-35.5,-143.5</position>
<gparam>LABEL_TEXT Y=A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>-71,-153.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>-74.5,-152.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>BA_NAND2</type>
<position>-51.5,-148.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>BA_NAND2</type>
<position>-62,-153.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>4.5,-97.5</position>
<gparam>LABEL_TEXT 4.NAND as NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>BA_NAND2</type>
<position>5,-105</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>-4,-105</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>38.5,-109.5</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>-7,-104</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>47,-109.5</position>
<gparam>LABEL_TEXT Y=A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>-4,-114.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>-7.5,-113.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>BA_NAND2</type>
<position>15.5,-109.5</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>BA_NAND2</type>
<position>5,-114.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>BA_NAND2</type>
<position>27.5,-109.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>47,-106.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>51,-106.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>5.5,-124.5</position>
<gparam>LABEL_TEXT 5.NAND as XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>BA_NAND2</type>
<position>29.5,-133.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>8.5,-132.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>51,-138</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>4.5,-132</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_TOGGLE</type>
<position>9,-144</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>BA_NAND2</type>
<position>40,-138</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>BA_NAND2</type>
<position>29.5,-143</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>BA_NAND2</type>
<position>18,-138</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>4.5,-143</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>60.5,-137.5</position>
<gparam>LABEL_TEXT Y=AB+BA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>58,-134.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>64.5,-134.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>9,-151.5</position>
<gparam>LABEL_TEXT 6.NAND as XNOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>BA_NAND2</type>
<position>20,-158</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_TOGGLE</type>
<position>-1,-157</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>185</ID>
<type>GA_LED</type>
<position>55,-162.5</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-5,-156.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-168.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>BA_NAND2</type>
<position>30.5,-162.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>BA_NAND2</type>
<position>20,-167.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>BA_NAND2</type>
<position>8.5,-162.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>-5,-167.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>68,-161.5</position>
<gparam>LABEL_TEXT Y=AB+BA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>72,-158</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>74.5,-158</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>BA_NAND2</type>
<position>42.5,-162.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>-3,-202</position>
<gparam>LABEL_TEXT NOR gate as a Universal gate</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>-56.5,-215.5</position>
<gparam>LABEL_TEXT 1.NOR gate as NOT gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_TOGGLE</type>
<position>-67,-224.5</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>206</ID>
<type>GA_LED</type>
<position>-47.5,-224.5</position>
<input>
<ID>N_in0</ID>109 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>-70,-224</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>-41.5,-224.5</position>
<gparam>LABEL_TEXT Y=A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>-39.5,-221.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>BE_NOR2</type>
<position>-57,-224.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>-57.5,-231</position>
<gparam>LABEL_TEXT 2.NOR gate as OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_TOGGLE</type>
<position>-67.5,-238</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_TOGGLE</type>
<position>-67.5,-244</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>-71.5,-237.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>-71.5,-243.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>BE_NOR2</type>
<position>-55.5,-240</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>BE_NOR2</type>
<position>-45.5,-240</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>GA_LED</type>
<position>-37,-240</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>-28,-239.5</position>
<gparam>LABEL_TEXT Y=A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>-56.5,-252</position>
<gparam>LABEL_TEXT 3.NOR gate as AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AA_TOGGLE</type>
<position>-67,-260</position>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_TOGGLE</type>
<position>-67,-268.5</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>-70.5,-259.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>-70.5,-268</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>BE_NOR2</type>
<position>-55,-260</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>BE_NOR2</type>
<position>-45,-263.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>GA_LED</type>
<position>-36,-263.5</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>-28,-262.5</position>
<gparam>LABEL_TEXT Y=A.B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>BE_NOR2</type>
<position>-55,-268.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>15,-214.5</position>
<gparam>LABEL_TEXT 4.NOR gate as NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>AA_TOGGLE</type>
<position>4.5,-222</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_TOGGLE</type>
<position>4.5,-230.5</position>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>1,-221.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>1,-230</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>BE_NOR2</type>
<position>16.5,-222</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>BE_NOR2</type>
<position>26.5,-225.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>GA_LED</type>
<position>45.5,-225.5</position>
<input>
<ID>N_in0</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>55,-225</position>
<gparam>LABEL_TEXT Y=A.B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>BE_NOR2</type>
<position>16.5,-230.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>BE_NOR2</type>
<position>36.5,-225.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_LABEL</type>
<position>55.5,-222</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>58.5,-222</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>14.5,-239</position>
<gparam>LABEL_TEXT 5.NOR gate as XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>4,-246</position>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>4,-256.5</position>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_LABEL</type>
<position>0.5,-246</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>1,-254</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>BE_NOR2</type>
<position>31,-247</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>BE_NOR2</type>
<position>41,-250.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>258</ID>
<type>GA_LED</type>
<position>60,-250.5</position>
<input>
<ID>N_in0</ID>141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>69.5,-250</position>
<gparam>LABEL_TEXT Y=AB+BA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>BE_NOR2</type>
<position>31,-255.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>261</ID>
<type>BE_NOR2</type>
<position>15.5,-250.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>67,-247</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>73.5,-247</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>BE_NOR2</type>
<position>50.5,-250.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>140 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>15.5,-263</position>
<gparam>LABEL_TEXT 6.NOR gate as XNOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_TOGGLE</type>
<position>0,-268.5</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_TOGGLE</type>
<position>0,-279</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>-3.5,-268.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>-3,-276.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>BE_NOR2</type>
<position>27,-269.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>BE_NOR2</type>
<position>37,-273</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>GA_LED</type>
<position>66.5,-273</position>
<input>
<ID>N_in0</ID>152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>AA_LABEL</type>
<position>80,-273</position>
<gparam>LABEL_TEXT Y=AB+BA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>BE_NOR2</type>
<position>27,-278</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>BE_NOR2</type>
<position>11.5,-273</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_LABEL</type>
<position>86,-270</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>AA_LABEL</type>
<position>84,-270</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>BE_NOR2</type>
<position>46.5,-273</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>BE_NOR2</type>
<position>57,-273</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_LABEL</type>
<position>-5.5,-297.5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>AA_TOGGLE</type>
<position>-75.5,-312</position>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>285</ID>
<type>AA_TOGGLE</type>
<position>-61.5,-312</position>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_LABEL</type>
<position>-68,-304.5</position>
<gparam>LABEL_TEXT 1.Using AOI gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_INVERTER</type>
<position>-70,-315.5</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_INVERTER</type>
<position>-57,-316.5</position>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>-75.5,-309</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>-61.5,-309</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND2</type>
<position>-35,-323</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND2</type>
<position>-34.5,-332.5</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_OR2</type>
<position>-24.5,-326.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>GA_LED</type>
<position>-17,-326.5</position>
<input>
<ID>N_in0</ID>159 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>AA_LABEL</type>
<position>-4.5,-325.5</position>
<gparam>LABEL_TEXT sum=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>AA_LABEL</type>
<position>-4.5,-322.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>AA_LABEL</type>
<position>4,-322.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>AA_AND2</type>
<position>-33.5,-341</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>GA_LED</type>
<position>-16.5,-340.5</position>
<input>
<ID>N_in0</ID>160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>AA_LABEL</type>
<position>-6.5,-340</position>
<gparam>LABEL_TEXT carry=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>30.5,-306</position>
<gparam>LABEL_TEXT 2.Using XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>AA_TOGGLE</type>
<position>17,-313.5</position>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_TOGGLE</type>
<position>31,-313.5</position>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>17,-310.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>AA_LABEL</type>
<position>31,-310.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>GA_LED</type>
<position>51.5,-321</position>
<input>
<ID>N_in2</ID>170 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>64,-320</position>
<gparam>LABEL_TEXT sum=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>AA_LABEL</type>
<position>64,-317</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>AA_LABEL</type>
<position>72.5,-316.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>43.5,-329.5</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>GA_LED</type>
<position>52.5,-329.5</position>
<input>
<ID>N_in0</ID>169 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>AA_LABEL</type>
<position>62.5,-329</position>
<gparam>LABEL_TEXT carry=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>331</ID>
<type>AI_XOR2</type>
<position>42,-321</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_LABEL</type>
<position>-64,-347.5</position>
<gparam>LABEL_TEXT 3.Using NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>333</ID>
<type>AA_TOGGLE</type>
<position>-75.5,-355.5</position>
<output>
<ID>OUT_0</ID>183 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_TOGGLE</type>
<position>-61.5,-355.5</position>
<output>
<ID>OUT_0</ID>185 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>340</ID>
<type>GA_LED</type>
<position>-26,-367</position>
<input>
<ID>N_in0</ID>191 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>341</ID>
<type>AA_LABEL</type>
<position>-14,-366</position>
<gparam>LABEL_TEXT sum=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>AA_LABEL</type>
<position>-14,-363</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>343</ID>
<type>AA_LABEL</type>
<position>-5.5,-363</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>345</ID>
<type>GA_LED</type>
<position>-24,-380.5</position>
<input>
<ID>N_in0</ID>193 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>AA_LABEL</type>
<position>-14,-380</position>
<gparam>LABEL_TEXT carry=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AA_LABEL</type>
<position>-75.5,-352.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>BA_NAND2</type>
<position>-56.5,-359.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_LABEL</type>
<position>-61.5,-352.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>BA_NAND2</type>
<position>-69,-360</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>BA_NAND2</type>
<position>-44,-364.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>BA_NAND2</type>
<position>-43.5,-371</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>BA_NAND2</type>
<position>-33.5,-367</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>BA_NAND2</type>
<position>-43,-380.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>BA_NAND2</type>
<position>-32.5,-380.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>35,-347.5</position>
<gparam>LABEL_TEXT 4.Using NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>AA_TOGGLE</type>
<position>21,-356.5</position>
<output>
<ID>OUT_0</ID>207 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_TOGGLE</type>
<position>38,-356.5</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>364</ID>
<type>GA_LED</type>
<position>80,-369.5</position>
<input>
<ID>N_in1</ID>217 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>88,-365.5</position>
<gparam>LABEL_TEXT sum=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>AA_LABEL</type>
<position>88,-362.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>367</ID>
<type>AA_LABEL</type>
<position>96,-362.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>GA_LED</type>
<position>72,-381.5</position>
<input>
<ID>N_in0</ID>218 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>369</ID>
<type>AA_LABEL</type>
<position>82.5,-381</position>
<gparam>LABEL_TEXT carry=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>AA_LABEL</type>
<position>20.5,-353.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>AA_LABEL</type>
<position>38,-353.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>BE_NOR2</type>
<position>27,-361.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>BE_NOR2</type>
<position>45,-360</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>BE_NOR2</type>
<position>55.5,-366</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>BE_NOR2</type>
<position>56,-374</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>BE_NOR2</type>
<position>65,-369.5</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>BE_NOR2</type>
<position>74,-369.5</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>386</ID>
<type>BE_NOR2</type>
<position>60.5,-381.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_LABEL</type>
<position>-31,-406</position>
<gparam>LABEL_TEXT HALF-SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,-380.5,-25,-380.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<connection>
<GID>345</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,-6,-50,-6</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-50,-7.5,-50,-6</points>
<intersection>-7.5 5</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-50,-7.5,-49,-7.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-50 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,-11,-50,-11</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>-50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-50,-11,-50,-9.5</points>
<intersection>-11 1</intersection>
<intersection>-9.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-50,-9.5,-49,-9.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-50 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-8.5,-39,-8.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-39 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-39,-8.5,-39,-8</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-373,21,-358.5</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<intersection>-373 3</intersection>
<intersection>-362.5 6</intersection>
<intersection>-360.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-360.5,24,-360.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21,-373,53,-373</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21,-362.5,24,-362.5</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-380.5,31,-361.5</points>
<intersection>-380.5 4</intersection>
<intersection>-365 2</intersection>
<intersection>-361.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-361.5,31,-361.5</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-365,52.5,-365</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>31,-380.5,57.5,-380.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-367,38,-358.5</points>
<connection>
<GID>363</GID>
<name>OUT_0</name></connection>
<intersection>-367 2</intersection>
<intersection>-361 3</intersection>
<intersection>-359 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38,-367,52.5,-367</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38,-361,42,-361</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38,-359,42,-359</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-382.5,50.5,-360</points>
<intersection>-382.5 4</intersection>
<intersection>-375 1</intersection>
<intersection>-360 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-375,53,-375</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-360,50.5,-360</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-382.5,57.5,-382.5</points>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-374,60.5,-370.5</points>
<intersection>-374 2</intersection>
<intersection>-370.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-370.5,62,-370.5</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-374,60.5,-374</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-368.5,60,-366</points>
<intersection>-368.5 1</intersection>
<intersection>-366 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-368.5,62,-368.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-366,60,-366</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-370.5,69.5,-368.5</points>
<intersection>-370.5 3</intersection>
<intersection>-369.5 2</intersection>
<intersection>-368.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-368.5,71,-368.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-369.5,69.5,-369.5</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>69.5,-370.5,71,-370.5</points>
<connection>
<GID>385</GID>
<name>IN_1</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-369.5,81,-369.5</points>
<connection>
<GID>364</GID>
<name>N_in1</name></connection>
<connection>
<GID>385</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63.5,-381.5,71,-381.5</points>
<connection>
<GID>386</GID>
<name>OUT</name></connection>
<connection>
<GID>368</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-101,-445.5,-101,-428</points>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection>
<intersection>-445.5 1</intersection>
<intersection>-429.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-101,-445.5,-63,-445.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>-101 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-101,-429.5,-98.5,-429.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-101 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,-456,-87,-428</points>
<connection>
<GID>390</GID>
<name>OUT_0</name></connection>
<intersection>-456 8</intersection>
<intersection>-438 1</intersection>
<intersection>-430.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,-438,-63.5,-438</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<intersection>-87 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-87,-430.5,-85.5,-430.5</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-87,-456,-61,-456</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-25,-52.5,-24</points>
<intersection>-25 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52.5,-25,-49,-25</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-56,-24,-52.5,-24</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92.5,-436,-63.5,-436</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>-92.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-92.5,-454,-92.5,-429.5</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>-454 7</intersection>
<intersection>-436 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-92.5,-454,-61,-454</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>-92.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-29,-52.5,-27</points>
<intersection>-29 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52.5,-27,-49,-27</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-56,-29,-52.5,-29</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79,-447.5,-79,-430.5</points>
<intersection>-447.5 2</intersection>
<intersection>-430.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-79.5,-430.5,-79,-430.5</points>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection>
<intersection>-79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,-447.5,-63,-447.5</points>
<connection>
<GID>397</GID>
<name>IN_1</name></connection>
<intersection>-79 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-439.5,-55,-437</points>
<intersection>-439.5 1</intersection>
<intersection>-437 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-439.5,-53,-439.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-437,-55,-437</points>
<connection>
<GID>396</GID>
<name>OUT</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-26,-38.5,-26</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-446.5,-55,-441.5</points>
<intersection>-446.5 2</intersection>
<intersection>-441.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-441.5,-53,-441.5</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-446.5,-55,-446.5</points>
<connection>
<GID>397</GID>
<name>OUT</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-440.5,-43.5,-440.5</points>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<connection>
<GID>399</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-435,-5,-429</points>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection>
<intersection>-435 6</intersection>
<intersection>-430.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-430.5,-1.5,-430.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-5,-435,23.5,-435</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection>
<intersection>-1.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-1.5,-435,-1.5,-432.5</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>-435 6</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-454,8.5,-429</points>
<connection>
<GID>411</GID>
<name>OUT_0</name></connection>
<intersection>-454 14</intersection>
<intersection>-443.5 3</intersection>
<intersection>-430 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-430,11,-430</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8.5,-443.5,24,-443.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>8.5 0</intersection>
<intersection>11 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>11,-443.5,11,-432</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>-443.5 3</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>8.5,-454,25,-454</points>
<connection>
<GID>427</GID>
<name>IN_1</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-437,17.5,-431</points>
<intersection>-437 1</intersection>
<intersection>-431 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-437,23.5,-437</points>
<connection>
<GID>422</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-431,17.5,-431</points>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56.5,-44.5,-48,-44.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-452,6,-431.5</points>
<intersection>-452 4</intersection>
<intersection>-441.5 1</intersection>
<intersection>-431.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-441.5,24,-441.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-431.5,6,-431.5</points>
<connection>
<GID>421</GID>
<name>OUT</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>6,-452,25,-452</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44,-44.5,-38,-44.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<connection>
<GID>93</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-437.5,31.5,-436</points>
<intersection>-437.5 1</intersection>
<intersection>-436 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-437.5,34,-437.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-436,31.5,-436</points>
<connection>
<GID>422</GID>
<name>OUT</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-69,-52,-68</points>
<intersection>-69 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-68,-47.5,-68</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-69,-52,-69</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-442.5,31.5,-439.5</points>
<intersection>-442.5 2</intersection>
<intersection>-439.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-439.5,34,-439.5</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-442.5,31.5,-442.5</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-66,-52,-64.5</points>
<intersection>-66 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-66,-47.5,-66</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-64.5,-52,-64.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-438.5,43.5,-438.5</points>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<connection>
<GID>412</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,-67,-38,-67</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<connection>
<GID>98</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-454,32.5,-452</points>
<intersection>-454 4</intersection>
<intersection>-453 1</intersection>
<intersection>-452 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-453,32.5,-453</points>
<connection>
<GID>427</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-452,34.5,-452</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>32.5,-454,34.5,-454</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-454,46,-453</points>
<connection>
<GID>416</GID>
<name>N_in2</name></connection>
<intersection>-453 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-453,46,-453</points>
<connection>
<GID>428</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-9,10.5,-8</points>
<intersection>-9 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-9,14.5,-9</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-8,10.5,-8</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-103.5,-500,-103.5,-477</points>
<connection>
<GID>431</GID>
<name>OUT_0</name></connection>
<intersection>-500 8</intersection>
<intersection>-491.5 3</intersection>
<intersection>-481 6</intersection>
<intersection>-479 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103.5,-479,-100.5,-479</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>-103.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-103.5,-491.5,-71.5,-491.5</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>-103.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-103.5,-481,-100.5,-481</points>
<connection>
<GID>441</GID>
<name>IN_1</name></connection>
<intersection>-103.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-103.5,-500,-71,-500</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>-103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-12.5,10.5,-11</points>
<intersection>-12.5 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-11,14.5,-11</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-12.5,10.5,-12.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-483.5,-93.5,-480</points>
<intersection>-483.5 2</intersection>
<intersection>-480 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-94.5,-480,-93.5,-480</points>
<connection>
<GID>441</GID>
<name>OUT</name></connection>
<intersection>-93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-93.5,-483.5,-72,-483.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-10,26.5,-9.5</points>
<connection>
<GID>104</GID>
<name>N_in3</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-10,26.5,-10</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,-485.5,-86.5,-477</points>
<connection>
<GID>432</GID>
<name>OUT_0</name></connection>
<intersection>-485.5 2</intersection>
<intersection>-479.5 3</intersection>
<intersection>-477.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,-485.5,-72,-485.5</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-86.5,-479.5,-82.5,-479.5</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-86.5,-477.5,-82.5,-477.5</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>-86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,-502,-74,-478.5</points>
<intersection>-502 6</intersection>
<intersection>-493.5 1</intersection>
<intersection>-478.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,-493.5,-71.5,-493.5</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>-74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76.5,-478.5,-74,-478.5</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<intersection>-74 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-74,-502,-71,-502</points>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>-74 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64,-492.5,-64,-489</points>
<intersection>-492.5 2</intersection>
<intersection>-489 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-489,-62.5,-489</points>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>-64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,-492.5,-64,-492.5</points>
<connection>
<GID>444</GID>
<name>OUT</name></connection>
<intersection>-64 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-487,-64.5,-484.5</points>
<intersection>-487 1</intersection>
<intersection>-484.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-487,-62.5,-487</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,-484.5,-64.5,-484.5</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-489,-55,-487</points>
<intersection>-489 3</intersection>
<intersection>-488 2</intersection>
<intersection>-487 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-487,-53.5,-487</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-56.5,-488,-55,-488</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55,-489,-53.5,-489</points>
<connection>
<GID>446</GID>
<name>IN_1</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-108.5,-65,-106.5</points>
<intersection>-108.5 2</intersection>
<intersection>-107.5 11</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-106.5,-63.5,-106.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65,-108.5,-63.5,-108.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-68,-107.5,-65,-107.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47.5,-488,-43.5,-488</points>
<connection>
<GID>446</GID>
<name>OUT</name></connection>
<connection>
<GID>433</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-108,-55,-107.5</points>
<intersection>-108 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-108,-52.5,-108</points>
<connection>
<GID>123</GID>
<name>N_in0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-107.5,-55,-107.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-65,-501,-50.5,-501</points>
<connection>
<GID>449</GID>
<name>OUT</name></connection>
<intersection>-50.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-50.5,-502,-50.5,-501</points>
<connection>
<GID>437</GID>
<name>N_in2</name></connection>
<intersection>-501 1</intersection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95,-606.5,-95,-535</points>
<connection>
<GID>452</GID>
<name>OUT_0</name></connection>
<intersection>-606.5 23</intersection>
<intersection>-598 14</intersection>
<intersection>-589.5 12</intersection>
<intersection>-568 6</intersection>
<intersection>-558.5 1</intersection>
<intersection>-536 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-95,-558.5,-51,-558.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>-95 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-95,-536,-93.5,-536</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>-95 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-95,-568,-50.5,-568</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>-95 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-95,-589.5,-49.5,-589.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-95 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-95,-598,-49.5,-598</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>-95 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-95,-606.5,-49.5,-606.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>-95 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-68,-123,-63.5,-123</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-63.5,-124,-63.5,-123</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-123 1</intersection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80.5,-608.5,-80.5,-535</points>
<connection>
<GID>453</GID>
<name>OUT_0</name></connection>
<intersection>-608.5 14</intersection>
<intersection>-600 10</intersection>
<intersection>-581.5 8</intersection>
<intersection>-570 6</intersection>
<intersection>-550.5 1</intersection>
<intersection>-536 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-80.5,-550.5,-51.5,-550.5</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-80.5,-536,-78,-536</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-80.5,-570,-50.5,-570</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-80.5,-581.5,-50,-581.5</points>
<connection>
<GID>481</GID>
<name>IN_1</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-80.5,-600,-49.5,-600</points>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-80.5,-608.5,-49.5,-608.5</points>
<connection>
<GID>495</GID>
<name>IN_1</name></connection>
<intersection>-80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,-127.5,-65.5,-126</points>
<intersection>-127.5 2</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,-126,-63.5,-126</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-67.5,-127.5,-65.5,-127.5</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-610.5,-64.5,-535.5</points>
<connection>
<GID>457</GID>
<name>OUT_0</name></connection>
<intersection>-610.5 14</intersection>
<intersection>-593.5 12</intersection>
<intersection>-583.5 8</intersection>
<intersection>-572 6</intersection>
<intersection>-542 1</intersection>
<intersection>-536.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-542,-52,-542</points>
<connection>
<GID>466</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-64.5,-536.5,-61.5,-536.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-64.5,-572,-50.5,-572</points>
<connection>
<GID>469</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-64.5,-583.5,-50,-583.5</points>
<connection>
<GID>481</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-64.5,-593.5,-49.5,-593.5</points>
<connection>
<GID>486</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-64.5,-610.5,-49.5,-610.5</points>
<connection>
<GID>495</GID>
<name>IN_2</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-538,-52,-538</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>-89.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-89.5,-579.5,-89.5,-536</points>
<connection>
<GID>462</GID>
<name>OUT_0</name></connection>
<intersection>-579.5 7</intersection>
<intersection>-548.5 5</intersection>
<intersection>-538 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-89.5,-548.5,-51.5,-548.5</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>-89.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-89.5,-579.5,-50,-579.5</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>-89.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-126,-55,-124</points>
<intersection>-126 2</intersection>
<intersection>-126 2</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-124,-53,-124</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-126,-53,-126</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>-57.5 3</intersection>
<intersection>-55 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-57.5,-126,-57.5,-125</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>-126 2</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73.5,-591.5,-73.5,-536</points>
<intersection>-591.5 6</intersection>
<intersection>-560.5 4</intersection>
<intersection>-540 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73.5,-540,-52,-540</points>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<intersection>-73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-74,-536,-73.5,-536</points>
<connection>
<GID>463</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-73.5,-560.5,-51,-560.5</points>
<connection>
<GID>468</GID>
<name>IN_1</name></connection>
<intersection>-73.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-73.5,-591.5,-49.5,-591.5</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>-73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-125,-43,-125</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<connection>
<GID>136</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-602,-56,-536.5</points>
<intersection>-602 6</intersection>
<intersection>-562.5 4</intersection>
<intersection>-552.5 1</intersection>
<intersection>-536.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-552.5,-51.5,-552.5</points>
<connection>
<GID>467</GID>
<name>IN_2</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-536.5,-56,-536.5</points>
<connection>
<GID>464</GID>
<name>OUT_0</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-56,-562.5,-51,-562.5</points>
<connection>
<GID>468</GID>
<name>IN_2</name></connection>
<intersection>-56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-56,-602,-49.5,-602</points>
<connection>
<GID>483</GID>
<name>IN_2</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,-550.5,-38.5,-547.5</points>
<intersection>-550.5 2</intersection>
<intersection>-547.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38.5,-547.5,-32,-547.5</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>-38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45.5,-550.5,-38.5,-550.5</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>-38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,-560.5,-38.5,-549.5</points>
<intersection>-560.5 2</intersection>
<intersection>-549.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38.5,-549.5,-32,-549.5</points>
<connection>
<GID>471</GID>
<name>IN_2</name></connection>
<intersection>-38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45,-560.5,-38.5,-560.5</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>-38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48.5,-148.5,-44.5,-148.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>-44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-44.5,-148.5,-44.5,-144</points>
<connection>
<GID>140</GID>
<name>N_in0</name></connection>
<intersection>-148.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,-570,-38.5,-551.5</points>
<intersection>-570 2</intersection>
<intersection>-551.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38.5,-551.5,-32,-551.5</points>
<connection>
<GID>471</GID>
<name>IN_3</name></connection>
<intersection>-38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-570,-38.5,-570</points>
<connection>
<GID>469</GID>
<name>OUT</name></connection>
<intersection>-38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-545.5,-39,-540</points>
<intersection>-545.5 1</intersection>
<intersection>-540 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-545.5,-32,-545.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>-39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46,-540,-39,-540</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25,-548.5,-18.5,-548.5</points>
<connection>
<GID>473</GID>
<name>N_in0</name></connection>
<connection>
<GID>471</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-585.5,-36,-581.5</points>
<intersection>-585.5 1</intersection>
<intersection>-581.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-585.5,-28,-585.5</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44,-581.5,-36,-581.5</points>
<connection>
<GID>481</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43.5,-587.5,-28,-587.5</points>
<connection>
<GID>488</GID>
<name>IN_1</name></connection>
<intersection>-43.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-43.5,-591.5,-43.5,-587.5</points>
<connection>
<GID>486</GID>
<name>OUT</name></connection>
<intersection>-587.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-154.5,-65,-152.5</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-153.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-153.5,-65,-153.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-600,-35.5,-589.5</points>
<intersection>-600 2</intersection>
<intersection>-589.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-589.5,-28,-589.5</points>
<connection>
<GID>488</GID>
<name>IN_2</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,-600,-35.5,-600</points>
<connection>
<GID>483</GID>
<name>OUT</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-145,-65,-143</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,-144,-65,-144</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-147.5,-56.5,-144</points>
<intersection>-147.5 1</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56.5,-147.5,-54.5,-147.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-59,-144,-56.5,-144</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,-588.5,-14.5,-587.5</points>
<connection>
<GID>489</GID>
<name>N_in3</name></connection>
<intersection>-588.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-588.5,-14.5,-588.5</points>
<connection>
<GID>488</GID>
<name>OUT</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-153.5,-56.5,-149.5</points>
<intersection>-153.5 2</intersection>
<intersection>-149.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56.5,-149.5,-54.5,-149.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-59,-153.5,-56.5,-153.5</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-608.5,-35.5,-591.5</points>
<intersection>-608.5 2</intersection>
<intersection>-591.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-591.5,-28,-591.5</points>
<connection>
<GID>488</GID>
<name>IN_3</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,-608.5,-35.5,-608.5</points>
<connection>
<GID>495</GID>
<name>OUT</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-115.5,2,-113.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,-114.5,2,-114.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-106,2,-104</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,-105,2,-105</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-108.5,10.5,-105</points>
<intersection>-108.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-108.5,12.5,-108.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-105,10.5,-105</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-114.5,10.5,-110.5</points>
<intersection>-114.5 2</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-110.5,12.5,-110.5</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-114.5,10.5,-114.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-110.5,24.5,-108.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-109.5,24.5,-109.5</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-109.5,37.5,-109.5</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<connection>
<GID>165</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-137,35,-133.5</points>
<intersection>-137 1</intersection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-137,37,-137</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-133.5,35,-133.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-143,35,-139</points>
<intersection>-143 2</intersection>
<intersection>-139 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-139,37,-139</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-143,35,-143</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-142,23.5,-134.5</points>
<intersection>-142 3</intersection>
<intersection>-138 2</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-134.5,26.5,-134.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-138,23.5,-138</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-142,26.5,-142</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-144,26.5,-144</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>15 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>15,-144,15,-139</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>-144 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-132.5,26.5,-132.5</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>15 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>15,-137,15,-132.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-132.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-138,50,-138</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<connection>
<GID>174</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-161.5,25.5,-158</points>
<intersection>-161.5 1</intersection>
<intersection>-158 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-161.5,27.5,-161.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-158,25.5,-158</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-167.5,25.5,-163.5</points>
<intersection>-167.5 2</intersection>
<intersection>-163.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-163.5,27.5,-163.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-167.5,25.5,-167.5</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-166.5,14,-159</points>
<intersection>-166.5 3</intersection>
<intersection>-162.5 2</intersection>
<intersection>-159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-159,17,-159</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-162.5,14,-162.5</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14,-166.5,17,-166.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-168.5,17,-168.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5.5,-168.5,5.5,-163.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>-168.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-157,17,-157</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>5.5 2</intersection>
<intersection>17 6</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>5.5,-161.5,5.5,-157</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-157 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>17,-157,17,-157</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-157 1</intersection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-163.5,39.5,-161.5</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-162.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-162.5,39.5,-162.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-162.5,54,-162.5</points>
<connection>
<GID>185</GID>
<name>N_in0</name></connection>
<connection>
<GID>195</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-225.5,-60,-223.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-224.5,-60,-224.5</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-224.5,-48.5,-224.5</points>
<connection>
<GID>206</GID>
<name>N_in0</name></connection>
<connection>
<GID>211</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-239,-62,-238</points>
<intersection>-239 1</intersection>
<intersection>-238 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-239,-58.5,-239</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,-238,-62,-238</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-244,-62,-241</points>
<intersection>-244 2</intersection>
<intersection>-241 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-241,-58.5,-241</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65.5,-244,-62,-244</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,-241,-48.5,-239</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-240 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52.5,-240,-48.5,-240</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>-48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42.5,-240,-38,-240</points>
<connection>
<GID>221</GID>
<name>N_in0</name></connection>
<connection>
<GID>220</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-261,-58,-259</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>-260 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-260,-58,-260</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-269.5,-58,-267.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-268.5,-58,-268.5</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,-262.5,-50,-260</points>
<intersection>-262.5 1</intersection>
<intersection>-260 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,-262.5,-48,-262.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-260,-50,-260</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>-50 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,-268.5,-50,-264.5</points>
<intersection>-268.5 2</intersection>
<intersection>-264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,-264.5,-48,-264.5</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>-50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-268.5,-50,-268.5</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>-50 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-263.5,-37,-263.5</points>
<connection>
<GID>230</GID>
<name>N_in0</name></connection>
<connection>
<GID>229</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-223,13.5,-221</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-222 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-222,13.5,-222</points>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-231.5,13.5,-229.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>-230.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-230.5,13.5,-230.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-224.5,21.5,-222</points>
<intersection>-224.5 1</intersection>
<intersection>-222 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-224.5,23.5,-224.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-222,21.5,-222</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-230.5,21.5,-226.5</points>
<intersection>-230.5 2</intersection>
<intersection>-226.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-226.5,23.5,-226.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-230.5,21.5,-230.5</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-226.5,33.5,-224.5</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-225.5,33.5,-225.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-225.5,44.5,-225.5</points>
<connection>
<GID>245</GID>
<name>N_in0</name></connection>
<connection>
<GID>248</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-249.5,36,-247</points>
<intersection>-249.5 1</intersection>
<intersection>-247 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-249.5,38,-249.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-247,36,-247</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-255.5,36,-251.5</points>
<intersection>-255.5 2</intersection>
<intersection>-251.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-251.5,38,-251.5</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-255.5,36,-255.5</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-246,28,-246</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12.5,-249.5,12.5,-246</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>-246 1</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-256.5,28,-256.5</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12.5,-256.5,12.5,-251.5</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>-256.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-254.5,23,-248</points>
<intersection>-254.5 3</intersection>
<intersection>-250.5 2</intersection>
<intersection>-248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-248,28,-248</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-250.5,23,-250.5</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23,-254.5,28,-254.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-251.5,47.5,-249.5</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>-250.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-250.5,47.5,-250.5</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-250.5,59,-250.5</points>
<connection>
<GID>258</GID>
<name>N_in0</name></connection>
<connection>
<GID>264</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-272,32,-269.5</points>
<intersection>-272 1</intersection>
<intersection>-269.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-272,34,-272</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-269.5,32,-269.5</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-278,32,-274</points>
<intersection>-278 2</intersection>
<intersection>-274 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-274,34,-274</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-278,32,-278</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-268.5,24,-268.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>8.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-272,8.5,-268.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>-268.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-279,24,-279</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>8.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8.5,-279,8.5,-274</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<intersection>-279 1</intersection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-277,19,-270.5</points>
<intersection>-277 3</intersection>
<intersection>-273 2</intersection>
<intersection>-270.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-270.5,24,-270.5</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-273,19,-273</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19,-277,24,-277</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-274,43.5,-272</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>-273 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-273,43.5,-273</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-274,54,-272</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>-273 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>49.5,-273,54,-273</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-273,65.5,-273</points>
<connection>
<GID>272</GID>
<name>N_in0</name></connection>
<connection>
<GID>279</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75.5,-340,-75.5,-314</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>-340 6</intersection>
<intersection>-331.5 1</intersection>
<intersection>-315.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75.5,-331.5,-37.5,-331.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-75.5,-315.5,-73,-315.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-75.5,-340,-36.5,-340</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-342,-61.5,-314</points>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>-342 6</intersection>
<intersection>-324 1</intersection>
<intersection>-316.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61.5,-324,-38,-324</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-61.5,-316.5,-60,-316.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-61.5,-342,-36.5,-342</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-67,-322,-38,-322</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>-67 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-67,-322,-67,-315.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>-322 1</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-333.5,-53.5,-316.5</points>
<intersection>-333.5 2</intersection>
<intersection>-316.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-316.5,-53.5,-316.5</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-333.5,-37.5,-333.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>-53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-325.5,-29.5,-323</points>
<intersection>-325.5 1</intersection>
<intersection>-323 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-325.5,-27.5,-325.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32,-323,-29.5,-323</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-332.5,-29.5,-327.5</points>
<intersection>-332.5 2</intersection>
<intersection>-327.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-327.5,-27.5,-327.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-31.5,-332.5,-29.5,-332.5</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21.5,-326.5,-18,-326.5</points>
<connection>
<GID>302</GID>
<name>N_in0</name></connection>
<connection>
<GID>300</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30.5,-341,-17.5,-341</points>
<connection>
<GID>309</GID>
<name>OUT</name></connection>
<intersection>-17.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-17.5,-341,-17.5,-340.5</points>
<connection>
<GID>311</GID>
<name>N_in0</name></connection>
<intersection>-341 1</intersection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-328.5,17,-315.5</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>-328.5 6</intersection>
<intersection>-320 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>17,-328.5,40.5,-328.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>17,-320,39,-320</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-330.5,31,-315.5</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>-330.5 6</intersection>
<intersection>-322 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>31,-330.5,40.5,-330.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31,-322,39,-322</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-329.5,51.5,-329.5</points>
<connection>
<GID>328</GID>
<name>N_in0</name></connection>
<connection>
<GID>327</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-322,51.5,-321</points>
<connection>
<GID>323</GID>
<name>N_in2</name></connection>
<intersection>-321 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-321,51.5,-321</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75.5,-379.5,-75.5,-357.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>-379.5 12</intersection>
<intersection>-363.5 6</intersection>
<intersection>-359 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75.5,-359,-72,-359</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-75.5,-363.5,-47,-363.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection>
<intersection>-72 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-72,-363.5,-72,-361</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>-363.5 6</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-75.5,-379.5,-46,-379.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>-75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-381.5,-61.5,-357.5</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>-381.5 11</intersection>
<intersection>-372 3</intersection>
<intersection>-358.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61.5,-358.5,-59.5,-358.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-61.5,-372,-46.5,-372</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>-61.5 0</intersection>
<intersection>-59.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-59.5,-372,-59.5,-360.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>-372 3</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-61.5,-381.5,-46,-381.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-365.5,-53,-359.5</points>
<intersection>-365.5 1</intersection>
<intersection>-359.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53,-365.5,-47,-365.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<intersection>-53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-359.5,-53,-359.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>-53 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-370,-64.5,-360</points>
<intersection>-370 1</intersection>
<intersection>-360 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,-370,-46.5,-370</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66,-360,-64.5,-360</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-366,-39,-364.5</points>
<intersection>-366 1</intersection>
<intersection>-364.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-366,-36.5,-366</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>-39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-41,-364.5,-39,-364.5</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-371,-39,-368</points>
<intersection>-371 2</intersection>
<intersection>-368 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-368,-36.5,-368</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>-39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-371,-39,-371</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30.5,-367,-27,-367</points>
<connection>
<GID>340</GID>
<name>N_in0</name></connection>
<connection>
<GID>357</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-381.5,-35.5,-379.5</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>-380.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,-380.5,-35.5,-380.5</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>